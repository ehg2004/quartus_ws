--library ieee;
--use ieee.std_logic_1164.all;
--
--package array_lab02_pkg is
--       	type array_4_bit_7 is array (6 downto 0) of std_logic_vector(3 downto 0);
--			type array_4_bit_6 is array (5 downto 0) of std_logic_vector(3 downto 0);
--		 -- type bus_array is array(natural range <>, natural range <>) of std_logic;
--end package;